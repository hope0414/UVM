import decode_in_pkg::*;
import decode_test_pkg::*;
import uvm_pkg::*;

module hvl_top;
  initial
  begin
 
    run_test("test_top");
  end
endmodule
