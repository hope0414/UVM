//----------------------------------------------------------------------
// Created with uvmf_gen version 2019.4_1
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// DESCRIPTION: 
// This file contains defines and typedefs to be compiled for use in
// the simulation running on the emulator when using Veloce.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
                                                                               

typedef logic [1:0] W_control_t;
typedef logic Mem_control_t;
typedef logic [5:0] E_control_t;
typedef logic [15:0] IR_t;
typedef logic [15:0] npc_out_t;

// pragma uvmf custom additional begin
// pragma uvmf custom additional end

