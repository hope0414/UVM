package decode_test_pkg;
  import uvm_pkg::*;
  //import questa_uvm_pkg::*;	
  import decode_in_pkg::*;

  `include "uvm_macros.svh"
  `include "test_top.sv"


endpackage
